`include "simple_mem.v"
`include "decoder_5to32.v"
`include "mux_4to1.v"
`include "mux_8to1.v"
`include "DFF.v"

module ram_32x32(clk,add_row,add_col,w_en,w_data,r_en,r_data);
   input clk,w_en,w_data,r_en;
   input [4:0] add_row,add_col;
   output      r_data;
   reg  data;
   wire [31:0]  row,colum;
   wire [31:0] 	d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31;
   wire [3:0] 	m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16,m17,m18,m19,m20,m21,m22,m23,m24,m25,m26,m27,m28,m29,m30,m31;
   wire [3:0] 	n;
   wire [31:0] 	sub_row,sub_colum;
   wire [4:0] 	address_row,address_col;
   wire 	write_en,read_en,write_data,read_data;

   
   decoder_5to32 ROW(add_row,sub_row);
   decoder_5to32 COL(add_col,sub_colum);

   DFF BUF00(clk,1'b0,w_en,write_en,);
   DFF BUF01(clk,1'b0,w_data,write_data,);
   DFF BUF10(clk,1'b0,r_en,read_en,);

   DFF BUF1[31:0] (clk,1'b0,sub_row[31:0],row[31:0],);
   DFF BUF2[31:0] (clk,1'b0,sub_colum[31:0],colum[31:0],);
   DFF BUF3[4:0] (clk,1'b0,add_row[4:0],address_row[4:0],);
   DFF BUF4[4:0] (clk,1'b0,add_col[4:0],address_col[4:0],);

   
   simple_mem MEM0[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0],row[0]}&colum[31:0],d0);
   
   simple_mem MEM1[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1],row[1]}&colum[31:0],d1);

   simple_mem MEM2[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2],row[2]}&colum[31:0],d2);
  
   simple_mem MEM3[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3],row[3]}&colum[31:0],d3);
   
   
   simple_mem MEM4[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4],row[4]}&colum[31:0],d4);
   
   simple_mem MEM5[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5],row[5]}&colum[31:0],d5);
   
   simple_mem MEM6[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6],row[6]}&colum[31:0],d6);
   
   simple_mem MEM7[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7],row[7]}&colum[31:0],d7);
   
   simple_mem MEM8[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8],row[8]}&colum[31:0],d8);
   
   simple_mem MEM9[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9],row[9]}&colum[31:0],d9);

   simple_mem MEM10[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10],row[10]}&colum[31:0],d10);
   
   simple_mem MEM11[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11],row[11]}&colum[31:0],d11);

   simple_mem MEM12[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12],row[12]}&colum[31:0],d12);
  
   simple_mem MEM13[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13],row[13]}&colum[31:0],d13);
   
   simple_mem MEM14[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14],row[14]}&colum[31:0],d14);
   
   simple_mem MEM15[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15],row[15]}&colum[31:0],d15);
   
   simple_mem MEM16[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16],row[16]}&colum[31:0],d16);
   
   simple_mem MEM17[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17],row[17]}&colum[31:0],d17);
   
   simple_mem MEM18[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18],row[18]}&colum[31:0],d18);
   
   simple_mem MEM19[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19],row[19]}&colum[31:0],d19);

   simple_mem MEM20[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20],row[20]}&colum[31:0],d20);
   
   simple_mem MEM21[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21],row[21]}&colum[31:0],d21);

   simple_mem MEM22[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22],row[22]}&colum[31:0],d22);
  
   simple_mem MEM23[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23],row[23]}&colum[31:0],d23);
   
   
   simple_mem MEM24[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24],row[24]}&colum[31:0],d24);
   
   simple_mem MEM25[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25],row[25]}&colum[31:0],d25);
   
   simple_mem MEM26[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26],row[26]}&colum[31:0],d26);
   
   simple_mem MEM27[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27],row[27]}&colum[31:0],d27);
   
   simple_mem MEM28[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28],row[28]}&colum[31:0],d28);
   
   simple_mem MEM29[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29],row[29]}&colum[31:0],d29);

   simple_mem MEM30[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30],row[30]}&colum[31:0],d30);
   
   simple_mem MEM31[31:0] (clk,{write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en,write_en}&{row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31]}&colum[31:0],write_data,{read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en,read_en}&{row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31],row[31]}&colum[31:0],d31);


   mux_8to1 MUX0(d0[0],d0[1],d0[2],d0[3],d0[4],d0[5],d0[6],d0[7],address_col[2:0],m0[0]);
   mux_8to1 MUX1(d0[8],d0[9],d0[10],d0[11],d0[12],d0[13],d0[14],d0[15],address_col[2:0],m0[1]);
   mux_8to1 MUX2(d0[16],d0[17],d0[18],d0[19],d0[20],d0[21],d0[22],d0[23],address_col[2:0],m0[2]);
   mux_8to1 MUX3(d0[24],d0[25],d0[26],d0[27],d0[28],d0[29],d0[30],d0[31],address_col[2:0],m0[3]);

   mux_4to1 MUX4(r0,m0[0],m0[1],m0[2],m0[3],address_col[4],address_col[3]);

   mux_8to1 MUX5(d1[0],d1[1],d1[2],d1[3],d1[4],d1[5],d1[6],d1[7],address_col[2:0],m1[0]);
   mux_8to1 MUX6(d1[8],d1[9],d1[10],d1[11],d1[12],d1[13],d1[14],d1[15],address_col[2:0],m1[1]);
   mux_8to1 MUX7(d1[16],d1[17],d1[18],d1[19],d1[20],d1[21],d1[22],d1[23],address_col[2:0],m1[2]);
   mux_8to1 MUX8(d1[24],d1[25],d1[26],d1[27],d1[28],d1[29],d1[30],d1[31],address_col[2:0],m1[3]);

   mux_4to1 MUX9(r1,m1[0],m1[1],m1[2],m1[3],address_col[4],address_col[3]);

   mux_8to1 MUX10(d2[0],d2[1],d2[2],d2[3],d2[4],d2[5],d2[6],d2[7],address_col[2:0],m2[0]);
   mux_8to1 MUX11(d2[8],d2[9],d2[10],d2[11],d2[12],d2[13],d2[14],d2[15],address_col[2:0],m2[1]);
   mux_8to1 MUX12(d2[16],d2[17],d2[18],d2[19],d2[20],d2[21],d2[22],d2[23],address_col[2:0],m2[2]);
   mux_8to1 MUX13(d2[24],d2[25],d2[26],d2[27],d2[28],d2[29],d2[30],d2[31],address_col[2:0],m2[3]);

   mux_4to1 MUX14(r2,m2[0],m2[1],m2[2],m2[3],address_col[4],address_col[3]);

   mux_8to1 MUX15(d3[0],d3[1],d3[2],d3[3],d3[4],d3[5],d3[6],d3[7],address_col[2:0],m3[0]);
   mux_8to1 MUX16(d3[8],d3[9],d3[10],d3[11],d3[12],d3[13],d3[14],d3[15],address_col[2:0],m3[1]);
   mux_8to1 MUX17(d3[16],d3[17],d3[18],d3[19],d3[20],d3[21],d3[22],d3[23],address_col[2:0],m3[2]);
   mux_8to1 MUX18(d3[24],d3[25],d3[26],d3[27],d3[28],d3[29],d3[30],d3[31],address_col[2:0],m3[3]);

   mux_4to1 MUX19(r3,m3[0],m3[1],m3[2],m3[3],address_col[4],address_col[3]);

   mux_8to1 MUX20(d4[0],d4[1],d4[2],d4[3],d4[4],d4[5],d4[6],d4[7],address_col[2:0],m4[0]);
   mux_8to1 MUX21(d4[8],d4[9],d4[10],d4[11],d4[12],d4[13],d4[14],d4[15],address_col[2:0],m4[1]);
   mux_8to1 MUX22(d4[16],d4[17],d4[18],d4[19],d4[20],d4[21],d4[22],d4[23],address_col[2:0],m4[2]);
   mux_8to1 MUX23(d4[24],d4[25],d4[26],d4[27],d4[28],d4[29],d4[30],d4[31],address_col[2:0],m4[3]);

   mux_4to1 MUX24(r4,m4[0],m4[1],m4[2],m4[3],address_col[4],address_col[3]);

   mux_8to1 MUX25(d5[0],d5[1],d5[2],d5[3],d5[4],d5[5],d5[6],d5[7],address_col[2:0],m5[0]);
   mux_8to1 MUX26(d5[8],d5[9],d5[10],d5[11],d5[12],d5[13],d5[14],d5[15],address_col[2:0],m5[1]);
   mux_8to1 MUX27(d5[16],d5[17],d5[18],d5[19],d5[20],d5[21],d5[22],d5[23],address_col[2:0],m5[2]);
   mux_8to1 MUX28(d5[24],d5[25],d5[26],d5[27],d5[28],d5[29],d5[30],d5[31],address_col[2:0],m5[3]);

   mux_4to1 MUX29(r5,m5[0],m5[1],m5[2],m5[3],address_col[4],address_col[3]);

   mux_8to1 MUX30(d6[0],d6[1],d6[2],d6[3],d6[4],d6[5],d6[6],d6[7],address_col[2:0],m6[0]);
   mux_8to1 MUX31(d6[8],d6[9],d6[10],d6[11],d6[12],d6[13],d6[14],d6[15],address_col[2:0],m6[1]);
   mux_8to1 MUX32(d6[16],d6[17],d6[18],d6[19],d6[20],d6[21],d6[22],d6[23],address_col[2:0],m6[2]);
   mux_8to1 MUX33(d6[24],d6[25],d6[26],d6[27],d6[28],d6[29],d6[30],d6[31],address_col[2:0],m6[3]);

   mux_4to1 MUX34(r6,m6[0],m6[1],m6[2],m6[3],address_col[4],address_col[3]);

   mux_8to1 MUX35(d7[0],d7[1],d7[2],d7[3],d7[4],d7[5],d7[6],d7[7],address_col[2:0],m7[0]);
   mux_8to1 MUX36(d7[8],d7[9],d7[10],d7[11],d7[12],d7[13],d7[14],d7[15],address_col[2:0],m7[1]);
   mux_8to1 MUX37(d7[16],d7[17],d7[18],d7[19],d7[20],d7[21],d7[22],d7[23],address_col[2:0],m7[2]);
   mux_8to1 MUX38(d7[24],d7[25],d7[26],d7[27],d7[28],d7[29],d7[30],d7[31],address_col[2:0],m7[3]);

   mux_4to1 MUX39(r7,m7[0],m7[1],m7[2],m7[3],address_col[4],address_col[3]);

   mux_8to1 MUX40(d8[0],d8[1],d8[2],d8[3],d8[4],d8[5],d8[6],d8[7],address_col[2:0],m8[0]);
   mux_8to1 MUX41(d8[8],d8[9],d8[10],d8[11],d8[12],d8[13],d8[14],d8[15],address_col[2:0],m8[1]);
   mux_8to1 MUX42(d8[16],d8[17],d8[18],d8[19],d8[20],d8[21],d8[22],d8[23],address_col[2:0],m8[2]);
   mux_8to1 MUX43(d8[24],d8[25],d8[26],d8[27],d8[28],d8[29],d8[30],d8[31],address_col[2:0],m8[3]);

   mux_4to1 MUX44(r8,m8[0],m8[1],m8[2],m8[3],address_col[4],address_col[3]);

   mux_8to1 MUX45(d9[0],d9[1],d9[2],d9[3],d9[4],d9[5],d9[6],d9[7],address_col[2:0],m9[0]);
   mux_8to1 MUX46(d9[8],d9[9],d9[10],d9[11],d9[12],d9[13],d9[14],d9[15],address_col[2:0],m9[1]);
   mux_8to1 MUX47(d9[16],d9[17],d9[18],d9[19],d9[20],d9[21],d9[22],d9[23],address_col[2:0],m9[2]);
   mux_8to1 MUX48(d9[24],d9[25],d9[26],d9[27],d9[28],d9[29],d9[30],d9[31],address_col[2:0],m9[3]);

   mux_4to1 MUX49(r9,m9[0],m9[1],m9[2],m9[3],address_col[4],address_col[3]);

   mux_8to1 MUX50(d10[0],d10[1],d10[2],d10[3],d10[4],d10[5],d10[6],d10[7],address_col[2:0],m10[0]);
   mux_8to1 MUX51(d10[8],d10[9],d10[10],d10[11],d10[12],d10[13],d10[14],d10[15],address_col[2:0],m10[1]);
   mux_8to1 MUX52(d10[16],d10[17],d10[18],d10[19],d10[20],d10[21],d10[22],d10[23],address_col[2:0],m10[2]);
   mux_8to1 MUX53(d10[24],d10[25],d10[26],d10[27],d10[28],d10[29],d10[30],d10[31],address_col[2:0],m10[3]);

   mux_4to1 MUX54(r10,m10[0],m10[1],m10[2],m10[3],address_col[4],address_col[3]);

   mux_8to1 MUX55(d11[0],d11[1],d11[2],d11[3],d11[4],d11[5],d11[6],d11[7],address_col[2:0],m11[0]);
   mux_8to1 MUX56(d11[8],d11[9],d11[10],d11[11],d11[12],d11[13],d11[14],d11[15],address_col[2:0],m11[1]);
   mux_8to1 MUX57(d11[16],d11[17],d11[18],d11[19],d11[20],d11[21],d11[22],d11[23],address_col[2:0],m11[2]);
   mux_8to1 MUX58(d11[24],d11[25],d11[26],d11[27],d11[28],d11[29],d11[30],d11[31],address_col[2:0],m11[3]);

   mux_4to1 MUX59(r11,m11[0],m11[1],m11[2],m11[3],address_col[4],address_col[3]);

   mux_8to1 MUX60(d12[0],d12[1],d12[2],d12[3],d12[4],d12[5],d12[6],d12[7],address_col[2:0],m12[0]);
   mux_8to1 MUX61(d12[8],d12[9],d12[10],d12[11],d12[12],d12[13],d12[14],d12[15],address_col[2:0],m12[1]);
   mux_8to1 MUX62(d12[16],d12[17],d12[18],d12[19],d12[20],d12[21],d12[22],d12[23],address_col[2:0],m12[2]);
   mux_8to1 MUX63(d12[24],d12[25],d12[26],d12[27],d12[28],d12[29],d12[30],d12[31],address_col[2:0],m12[3]);

   mux_4to1 MUX64(r12,m12[0],m12[1],m12[2],m12[3],address_col[4],address_col[3]);

   mux_8to1 MUX65(d13[0],d13[1],d13[2],d13[3],d13[4],d13[5],d13[6],d13[7],address_col[2:0],m13[0]);
   mux_8to1 MUX66(d13[8],d13[9],d13[10],d13[11],d13[12],d13[13],d13[14],d13[15],address_col[2:0],m13[1]);
   mux_8to1 MUX67(d13[16],d13[17],d13[18],d13[19],d13[20],d13[21],d13[22],d13[23],address_col[2:0],m13[2]);
   mux_8to1 MUX68(d13[24],d13[25],d13[26],d13[27],d13[28],d13[29],d13[30],d13[31],address_col[2:0],m13[3]);

   mux_4to1 MUX69(r13,m13[0],m13[1],m13[2],m13[3],address_col[4],address_col[3]);

   mux_8to1 MUX70(d14[0],d14[1],d14[2],d14[3],d14[4],d14[5],d14[6],d14[7],address_col[2:0],m14[0]);
   mux_8to1 MUX71(d14[8],d14[9],d14[10],d14[11],d14[12],d14[13],d14[14],d14[15],address_col[2:0],m14[1]);
   mux_8to1 MUX72(d14[16],d14[17],d14[18],d14[19],d14[20],d14[21],d14[22],d14[23],address_col[2:0],m14[2]);
   mux_8to1 MUX73(d14[24],d14[25],d14[26],d14[27],d14[28],d14[29],d14[30],d14[31],address_col[2:0],m14[3]);

   mux_4to1 MUX74(r14,m14[0],m14[1],m14[2],m14[3],address_col[4],address_col[3]);

   mux_8to1 MUX75(d15[0],d15[1],d15[2],d15[3],d15[4],d15[5],d15[6],d15[7],address_col[2:0],m15[0]);
   mux_8to1 MUX76(d15[8],d15[9],d15[10],d15[11],d15[12],d15[13],d15[14],d15[15],address_col[2:0],m15[1]);
   mux_8to1 MUX77(d15[16],d15[17],d15[18],d15[19],d15[20],d15[21],d15[22],d15[23],address_col[2:0],m15[2]);
   mux_8to1 MUX78(d15[24],d15[25],d15[26],d15[27],d15[28],d15[29],d15[30],d15[31],address_col[2:0],m15[3]);

   mux_4to1 MUX79(r15,m15[0],m15[1],m15[2],m15[3],address_col[4],address_col[3]);

   mux_8to1 MUX80(d16[0],d16[1],d16[2],d16[3],d16[4],d16[5],d16[6],d16[7],address_col[2:0],m16[0]);
   mux_8to1 MUX81(d16[8],d16[9],d16[10],d16[11],d16[12],d16[13],d16[14],d16[15],address_col[2:0],m16[1]);
   mux_8to1 MUX82(d16[16],d16[17],d16[18],d16[19],d16[20],d16[21],d16[22],d16[23],address_col[2:0],m16[2]);
   mux_8to1 MUX83(d16[24],d16[25],d16[26],d16[27],d16[28],d16[29],d16[30],d16[31],address_col[2:0],m16[3]);

   mux_4to1 MUX84(r16,m16[0],m16[1],m16[2],m16[3],address_col[4],address_col[3]);

   mux_8to1 MUX85(d17[0],d17[1],d17[2],d17[3],d17[4],d17[5],d17[6],d17[7],address_col[2:0],m17[0]);
   mux_8to1 MUX86(d17[8],d17[9],d17[10],d17[11],d17[12],d17[13],d17[14],d17[15],address_col[2:0],m17[1]);
   mux_8to1 MUX87(d17[16],d17[17],d17[18],d17[19],d17[20],d17[21],d17[22],d17[23],address_col[2:0],m17[2]);
   mux_8to1 MUX88(d17[24],d17[25],d17[26],d17[27],d17[28],d17[29],d17[30],d17[31],address_col[2:0],m17[3]);

   mux_4to1 MUX89(r17,m17[0],m17[1],m17[2],m17[3],address_col[4],address_col[3]);

   mux_8to1 MUX90(d18[0],d18[1],d18[2],d18[3],d18[4],d18[5],d18[6],d18[7],address_col[2:0],m18[0]);
   mux_8to1 MUX91(d18[8],d18[9],d18[10],d18[11],d18[12],d18[13],d18[14],d18[15],address_col[2:0],m18[1]);
   mux_8to1 MUX92(d18[16],d18[17],d18[18],d18[19],d18[20],d18[21],d18[22],d18[23],address_col[2:0],m18[2]);
   mux_8to1 MUX93(d18[24],d18[25],d18[26],d18[27],d18[28],d18[29],d18[30],d18[31],address_col[2:0],m18[3]);

   mux_4to1 MUX94(r18,m18[0],m18[1],m18[2],m18[3],address_col[4],address_col[3]);

   mux_8to1 MUX95(d19[0],d19[1],d19[2],d19[3],d19[4],d19[5],d19[6],d19[7],address_col[2:0],m19[0]);
   mux_8to1 MUX96(d19[8],d19[9],d19[10],d19[11],d19[12],d19[13],d19[14],d19[15],address_col[2:0],m19[1]);
   mux_8to1 MUX97(d19[16],d19[17],d19[18],d19[19],d19[20],d19[21],d19[22],d19[23],address_col[2:0],m19[2]);
   mux_8to1 MUX98(d19[24],d19[25],d19[26],d19[27],d19[28],d19[29],d19[30],d19[31],address_col[2:0],m19[3]);

   mux_4to1 MUX99(r19,m19[0],m19[1],m19[2],m19[3],address_col[4],address_col[3]);

   mux_8to1 MUX100(d20[0],d20[1],d20[2],d20[3],d20[4],d20[5],d20[6],d20[7],address_col[2:0],m20[0]);
   mux_8to1 MUX101(d20[8],d20[9],d20[10],d20[11],d20[12],d20[13],d20[14],d20[15],address_col[2:0],m20[1]);
   mux_8to1 MUX102(d20[16],d20[17],d20[18],d20[19],d20[20],d20[21],d20[22],d20[23],address_col[2:0],m20[2]);
   mux_8to1 MUX103(d20[24],d20[25],d20[26],d20[27],d20[28],d20[29],d20[30],d20[31],address_col[2:0],m20[3]);

   mux_4to1 MUX104(r20,m20[0],m20[1],m20[2],m20[3],address_col[4],address_col[3]);

   mux_8to1 MUX105(d21[0],d21[1],d21[2],d21[3],d21[4],d21[5],d21[6],d21[7],address_col[2:0],m21[0]);
   mux_8to1 MUX106(d21[8],d21[9],d21[10],d21[11],d21[12],d21[13],d21[14],d21[15],address_col[2:0],m21[1]);
   mux_8to1 MUX107(d21[16],d21[17],d21[18],d21[19],d21[20],d21[21],d21[22],d21[23],address_col[2:0],m21[2]);
   mux_8to1 MUX108(d21[24],d21[25],d21[26],d21[27],d21[28],d21[29],d21[30],d21[31],address_col[2:0],m21[3]);

   mux_4to1 MUX109(r21,m21[0],m21[1],m21[2],m21[3],address_col[4],address_col[3]);

   mux_8to1 MUX110(d22[0],d22[1],d22[2],d22[3],d22[4],d22[5],d22[6],d22[7],address_col[2:0],m22[0]);
   mux_8to1 MUX111(d22[8],d22[9],d22[10],d22[11],d22[12],d22[13],d22[14],d22[15],address_col[2:0],m22[1]);
   mux_8to1 MUX112(d22[16],d22[17],d22[18],d22[19],d22[20],d22[21],d22[22],d22[23],address_col[2:0],m22[2]);
   mux_8to1 MUX113(d22[24],d22[25],d22[26],d22[27],d22[28],d22[29],d22[30],d22[31],address_col[2:0],m22[3]);

   mux_4to1 MUX114(r22,m22[0],m22[1],m22[2],m22[3],address_col[4],address_col[3]);

   mux_8to1 MUX115(d23[0],d23[1],d23[2],d23[3],d23[4],d23[5],d23[6],d23[7],address_col[2:0],m23[0]);
   mux_8to1 MUX116(d23[8],d23[9],d23[10],d23[11],d23[12],d23[13],d23[14],d23[15],address_col[2:0],m23[1]);
   mux_8to1 MUX117(d23[16],d23[17],d23[18],d23[19],d23[20],d23[21],d23[22],d23[23],address_col[2:0],m23[2]);
   mux_8to1 MUX118(d23[24],d23[25],d23[26],d23[27],d23[28],d23[29],d23[30],d23[31],address_col[2:0],m23[3]);

   mux_4to1 MUX119(r23,m23[0],m23[1],m23[2],m23[3],address_col[4],address_col[3]);

   mux_8to1 MUX120(d24[0],d24[1],d24[2],d24[3],d24[4],d24[5],d24[6],d24[7],address_col[2:0],m24[0]);
   mux_8to1 MUX121(d24[8],d24[9],d24[10],d24[11],d24[12],d24[13],d24[14],d24[15],address_col[2:0],m24[1]);
   mux_8to1 MUX122(d24[16],d24[17],d24[18],d24[19],d24[20],d24[21],d24[22],d24[23],address_col[2:0],m24[2]);
   mux_8to1 MUX123(d24[24],d24[25],d24[26],d24[27],d24[28],d24[29],d24[30],d24[31],address_col[2:0],m24[3]);

   mux_4to1 MUX124(r24,m24[0],m24[1],m24[2],m24[3],address_col[4],address_col[3]);

   mux_8to1 MUX125(d25[0],d25[1],d25[2],d25[3],d25[4],d25[5],d25[6],d25[7],address_col[2:0],m25[0]);
   mux_8to1 MUX126(d25[8],d25[9],d25[10],d25[11],d25[12],d25[13],d25[14],d25[15],address_col[2:0],m25[1]);
   mux_8to1 MUX127(d25[16],d25[17],d25[18],d25[19],d25[20],d25[21],d25[22],d25[23],address_col[2:0],m25[2]);
   mux_8to1 MUX128(d25[24],d25[25],d25[26],d25[27],d25[28],d25[29],d25[30],d25[31],address_col[2:0],m25[3]);

   mux_4to1 MUX129(r25,m25[0],m25[1],m25[2],m25[3],address_col[4],address_col[3]);

   mux_8to1 MUX130(d26[0],d26[1],d26[2],d26[3],d26[4],d26[5],d26[6],d26[7],address_col[2:0],m26[0]);
   mux_8to1 MUX131(d26[8],d26[9],d26[10],d26[11],d26[12],d26[13],d26[14],d26[15],address_col[2:0],m26[1]);
   mux_8to1 MUX132(d26[16],d26[17],d26[18],d26[19],d26[20],d26[21],d26[22],d26[23],address_col[2:0],m26[2]);
   mux_8to1 MUX133(d26[24],d26[25],d26[26],d26[27],d26[28],d26[29],d26[30],d26[31],address_col[2:0],m26[3]);

   mux_4to1 MUX134(r26,m26[0],m26[1],m26[2],m26[3],address_col[4],address_col[3]);

   mux_8to1 MUX135(d27[0],d27[1],d27[2],d27[3],d27[4],d27[5],d27[6],d27[7],address_col[2:0],m27[0]);
   mux_8to1 MUX136(d27[8],d27[9],d27[10],d27[11],d27[12],d27[13],d27[14],d27[15],address_col[2:0],m27[1]);
   mux_8to1 MUX137(d27[16],d27[17],d27[18],d27[19],d27[20],d27[21],d27[22],d27[23],address_col[2:0],m27[2]);
   mux_8to1 MUX138(d27[24],d27[25],d27[26],d27[27],d27[28],d27[29],d27[30],d27[31],address_col[2:0],m27[3]);

   mux_4to1 MUX139(r27,m27[0],m27[1],m27[2],m27[3],address_col[4],address_col[3]);

   mux_8to1 MUX140(d28[0],d28[1],d28[2],d28[3],d28[4],d28[5],d28[6],d28[7],address_col[2:0],m28[0]);
   mux_8to1 MUX141(d28[8],d28[9],d28[10],d28[11],d28[12],d28[13],d28[14],d28[15],address_col[2:0],m28[1]);
   mux_8to1 MUX142(d28[16],d28[17],d28[18],d28[19],d28[20],d28[21],d28[22],d28[23],address_col[2:0],m28[2]);
   mux_8to1 MUX143(d28[24],d28[25],d28[26],d28[27],d28[28],d28[29],d28[30],d28[31],address_col[2:0],m28[3]);

   mux_4to1 MUX144(r28,m28[0],m28[1],m28[2],m28[3],address_col[4],address_col[3]);

   mux_8to1 MUX145(d29[0],d29[1],d29[2],d29[3],d29[4],d29[5],d29[6],d29[7],address_col[2:0],m29[0]);
   mux_8to1 MUX146(d29[8],d29[9],d29[10],d29[11],d29[12],d29[13],d29[14],d29[15],address_col[2:0],m29[1]);
   mux_8to1 MUX147(d29[16],d29[17],d29[18],d29[19],d29[20],d29[21],d29[22],d29[23],address_col[2:0],m29[2]);
   mux_8to1 MUX148(d29[24],d29[25],d29[26],d29[27],d29[28],d29[29],d29[30],d29[31],address_col[2:0],m29[3]);

   mux_4to1 MUX149(r29,m29[0],m29[1],m29[2],m29[3],address_col[4],address_col[3]);


   mux_8to1 MUX150(d30[0],d30[1],d30[2],d30[3],d30[4],d30[5],d30[6],d30[7],address_col[2:0],m30[0]);
   mux_8to1 MUX151(d30[8],d30[9],d30[10],d30[11],d30[12],d30[13],d30[14],d30[15],address_col[2:0],m30[1]);
   mux_8to1 MUX152(d30[16],d30[17],d30[18],d30[19],d30[20],d30[21],d30[22],d30[23],address_col[2:0],m30[2]);
   mux_8to1 MUX153(d30[24],d30[25],d30[26],d30[27],d30[28],d30[29],d30[30],d30[31],address_col[2:0],m30[3]);

   mux_4to1 MUX154(r30,m30[0],m30[1],m30[2],m30[3],address_col[4],address_col[3]);

   mux_8to1 MUX155(d31[0],d31[1],d31[2],d31[3],d31[4],d31[5],d31[6],d31[7],address_col[2:0],m31[0]);
   mux_8to1 MUX156(d31[8],d31[9],d31[10],d31[11],d31[12],d31[13],d31[14],d31[15],address_col[2:0],m31[1]);
   mux_8to1 MUX157(d31[16],d31[17],d31[18],d31[19],d31[20],d31[21],d31[22],d31[23],address_col[2:0],m31[2]);
   mux_8to1 MUX158(d31[24],d31[25],d31[26],d31[27],d31[28],d31[29],d31[30],d31[31],address_col[2:0],m31[3]);

   mux_4to1 MUX159(r31,m31[0],m31[1],m31[2],m31[3],address_col[4],address_col[3]);
   



   mux_8to1 MUX160(r0,r1,r2,r3,r4,r5,r6,r7,address_row[2:0],n[0]);
   mux_8to1 MUX161(r8,r9,r10,r11,r12,r13,r14,r15,address_row[2:0],n[1]);
   mux_8to1 MUX162(r16,r17,r18,r19,r20,r21,r22,r23,address_row[2:0],n[2]);
   mux_8to1 MUX163(r24,r25,r26,r27,r28,r29,r30,r31,address_row[2:0],n[3]);

   mux_4to1 MUX164(r_data,n[0],n[1],n[2],n[3],address_row[4],address_row[3]);


endmodule // ram_32x32

   
